library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Correlation_Gate is
	generic(
	input_size : integer := 0
	);
	port(
		CLK : in std_logic := '0';
		input_func : in std_logic_vector(input_size*8-1 downto 0) := (others => '0');
		input_adc : in std_logic_vector(input_Size*8-1 downto 0) := (others => '0');
		output : out std_logic_vector(18 downto 0) := (others => '0')
	);
end entity;

architecture arc of Correlation_Gate is

begin

process(CLK)
variable o : integer range 0 to 300000 := 0;
begin
	if(rising_edge(CLK)) then
		o := 0;
		for i in 1 to input_size loop
			o := o + (to_integer(unsigned((input_adc(i*8-1 downto i*8-8)))) * to_integer(unsigned((input_func(i*8-1 downto i*8-8)))));
		end loop;
		output <= std_logic_vector(to_unsigned(o, output'length));
	end if;
end process;

end architecture;