-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.0.1 Build 232 06/12/2013 Service Pack 1 SJ Web Edition
-- Created on Thu Jan 05 12:46:30 2023

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY StateMachineWizard IS
    PORT (
        reset : IN STD_LOGIC := '0';
        clock : IN STD_LOGIC;
        doneReadMemory : IN STD_LOGIC := '0';
        start : IN STD_LOGIC := '0';
        readMemoryEN : OUT STD_LOGIC;
        searchSignalEN : OUT STD_LOGIC
    );
END StateMachineWizard;

ARCHITECTURE BEHAVIOR OF StateMachineWizard IS
    TYPE type_fstate IS (idleState,readMemoryState,readSignalState);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,doneReadMemory,start)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= idleState;
            readMemoryEN <= '0';
            searchSignalEN <= '0';
        ELSE
            readMemoryEN <= '0';
            searchSignalEN <= '0';
            CASE fstate IS
                WHEN idleState =>
                    IF ((start = '1')) THEN
                        reg_fstate <= readMemoryState;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= idleState;
                    END IF;
                WHEN readMemoryState =>
                    IF ((doneReadMemory = '1')) THEN
                        reg_fstate <= readSignalState;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= readMemoryState;
                    END IF;

                    readMemoryEN <= '1';
                WHEN readSignalState =>
                    IF ((start = '0')) THEN
                        reg_fstate <= idleState;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= readSignalState;
                    END IF;

                    searchSignalEN <= '1';
                WHEN OTHERS => 
                    readMemoryEN <= 'X';
                    searchSignalEN <= 'X';
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
